`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: ICT 
// 
// Create Date: 20:54:07 05/07/2015 
// Design Name: Multiple constant rotations design
// Module Name: main 
// Project Name: MCR - Multiplierless  Constant Rotators Based on Combined Coefficient Selection and Shift and add Implementation
// Target Devices: FPGA Spartan 3E-500 nexys 2
// Description: 
//			This code implements Multiple constant rotation design. It takes 2 angles, R_fixed,maximum usable number of adders and 
//			maximum allowable error as input and gives optimum most coordinates of specified angle with respect to origin.
//////////////////////////////////////////////////////////////////////////////////

module main(clk,R_fixed,angle1,adder,error,angle2,final_cord1,final_cord2
    );
	
wire [13:0] R_LUT[255:0];
wire [13:0] tan_LUT[255:0];
wire [3:0] adder_LUT[255:0];
wire [13:0] sind_LUT[19:0];

/*****************************************************************/
//Error Index Look up table
assign sind_LUT[0]=14'b00000001001001;
assign sind_LUT[1]=14'b00000001010000;
assign sind_LUT[2]=14'b00000001011000;
assign sind_LUT[3]=14'b00000001011111;
assign sind_LUT[4]=14'b00000001100110;
assign sind_LUT[5]=14'b00000001101110;
assign sind_LUT[6]=14'b00000001110101;
assign sind_LUT[7]=14'b00000001111100;
assign sind_LUT[8]=14'b00000010000100;
assign sind_LUT[9]=14'b00000010001011;
assign sind_LUT[10]=14'b00000010010010;
assign sind_LUT[11]=14'b00000010011010;
assign sind_LUT[12]=14'b00000010100001;
assign sind_LUT[13]=14'b00000010101000;
assign sind_LUT[14]=14'b00000010110000;
assign sind_LUT[15]=14'b00000010110111;
assign sind_LUT[16]=14'b00000010111110;
assign sind_LUT[17]=14'b00000011000110;
assign sind_LUT[18]=14'b00000011001101;
assign sind_LUT[19]=14'b00000011010100;

/*****************************************************************/
//R Look up table
assign R_LUT[0]=14'b000000000000000;
assign R_LUT[1]=14'b000000010000000;
assign R_LUT[2]=14'b000000100000000;
assign R_LUT[3]=14'b000000110000000;
assign R_LUT[4]=14'b000001000000000;
assign R_LUT[5]=14'b000001010000000;
assign R_LUT[6]=14'b000001100000000;
assign R_LUT[7]=14'b000001110000000;
assign R_LUT[8]=14'b000010000000000;
assign R_LUT[9]=14'b000010010000000;
assign R_LUT[10]=14'b00010100000000;
assign R_LUT[11]=14'b00010110000000;
assign R_LUT[12]=14'b00011000000000;
assign R_LUT[13]=14'b00011010000000;
assign R_LUT[14]=14'b00011100000000;
assign R_LUT[15]=14'b00011110000000;
assign R_LUT[16]=14'b00000010000000;
assign R_LUT[17]=14'b00000010110101;
assign R_LUT[18]=14'b00000100011110;
assign R_LUT[19]=14'b00000110010100;
assign R_LUT[20]=14'b00001000001111;
assign R_LUT[21]=14'b00001010001100;
assign R_LUT[22]=14'b00001100001010;
assign R_LUT[23]=14'b00001110001001;
assign R_LUT[24]=14'b00010000000111;
assign R_LUT[25]=14'b00010010000111;
assign R_LUT[26]=14'b00010100000110;
assign R_LUT[27]=14'b00010110000101;
assign R_LUT[28]=14'b00011000000101;
assign R_LUT[29]=14'b00011010000100;
assign R_LUT[30]=14'b00011100000100;
assign R_LUT[31]=14'b00011110000100;
assign R_LUT[32]=14'b00000100000000;
assign R_LUT[33]=14'b00000100011110;
assign R_LUT[34]=14'b00000101101010;
assign R_LUT[35]=14'b00000111001101;
assign R_LUT[36]=14'b00001000111100;
assign R_LUT[37]=14'b00001010110001;
assign R_LUT[38]=14'b00001100101001;
assign R_LUT[39]=14'b00001110100011;
assign R_LUT[40]=14'b00010000011111;
assign R_LUT[41]=14'b00010010011100;
assign R_LUT[42]=14'b00010100011001;
assign R_LUT[43]=14'b00010110010111;
assign R_LUT[44]=14'b00011000010101;
assign R_LUT[45]=14'b00011010010011;
assign R_LUT[46]=14'b00011100010010;
assign R_LUT[47]=14'b00011110010000;
assign R_LUT[48]=14'b00000110000000;
assign R_LUT[49]=14'b00000110010100;
assign R_LUT[50]=14'b00000111001101;
assign R_LUT[51]=14'b00001000011111;
assign R_LUT[52]=14'b00001010000000;
assign R_LUT[53]=14'b00001011101010;
assign R_LUT[54]=14'b00001101011010;
assign R_LUT[55]=14'b00001111001110;
assign R_LUT[56]=14'b00010001000101;
assign R_LUT[57]=14'b00010010111110;
assign R_LUT[58]=14'b00010100111000;
assign R_LUT[59]=14'b00010110110011;
assign R_LUT[60]=14'b00011000101111;
assign R_LUT[61]=14'b00011010101011;
assign R_LUT[62]=14'b00011100101000;
assign R_LUT[63]=14'b00011110100110;
assign R_LUT[64]=14'b00001000000000;
assign R_LUT[65]=14'b00001000001111;
assign R_LUT[66]=14'b00001000111100;
assign R_LUT[67]=14'b00001010000000;
assign R_LUT[68]=14'b00001011010100;
assign R_LUT[69]=14'b00001100110011;
assign R_LUT[70]=14'b00001110011011;
assign R_LUT[71]=14'b00010000000111;
assign R_LUT[72]=14'b00010001111000;
assign R_LUT[73]=14'b00010011101100;
assign R_LUT[74]=14'b00010101100010;
assign R_LUT[75]=14'b00010111011010;
assign R_LUT[76]=14'b00011001010011;
assign R_LUT[77]=14'b00011011001100;
assign R_LUT[78]=14'b00011101000111;
assign R_LUT[79]=14'b00011111000011;
assign R_LUT[80]=14'b00001010000000;
assign R_LUT[81]=14'b00001010001100;
assign R_LUT[82]=14'b00001010110001;
assign R_LUT[83]=14'b00001011101010;
assign R_LUT[84]=14'b00001100110011;
assign R_LUT[85]=14'b00001110001001;
assign R_LUT[86]=14'b00001111100111;
assign R_LUT[87]=14'b00010001001101;
assign R_LUT[88]=14'b00010010110111;
assign R_LUT[89]=14'b00010100100101;
assign R_LUT[90]=14'b00010110010111;
assign R_LUT[91]=14'b00011000001010;
assign R_LUT[92]=14'b00011010000000;
assign R_LUT[93]=14'b00011011110110;
assign R_LUT[94]=14'b00011101101110;
assign R_LUT[95]=14'b00011111100111;
assign R_LUT[96]=14'b00001100000000;
assign R_LUT[97]=14'b00001100001010;
assign R_LUT[98]=14'b00001100101001;
assign R_LUT[99]=14'b00001101011010;
assign R_LUT[100]=14'b00001110011011;
assign R_LUT[101]=14'b00001111100111;
assign R_LUT[102]=14'b00010000111110;
assign R_LUT[103]=14'b00010010011100;
assign R_LUT[104]=14'b00010100000000;
assign R_LUT[105]=14'b00010101101000;
assign R_LUT[106]=14'b00010111010100;
assign R_LUT[107]=14'b00011001000011;
assign R_LUT[108]=14'b00011010110101;
assign R_LUT[109]=14'b00011100101000;
assign R_LUT[110]=14'b00011110011101;
assign R_LUT[111]=14'b00100000010011;
assign R_LUT[112]=14'b00001110000000;
assign R_LUT[113]=14'b00001110001001;
assign R_LUT[114]=14'b00001110100011;
assign R_LUT[115]=14'b00001111001110;
assign R_LUT[116]=14'b00010000000111;
assign R_LUT[117]=14'b00010001001101;
assign R_LUT[118]=14'b00010010011100;
assign R_LUT[119]=14'b00010011110011;
assign R_LUT[120]=14'b00010101010000;
assign R_LUT[121]=14'b00010110110011;
assign R_LUT[122]=14'b00011000011010;
assign R_LUT[123]=14'b00011010000100;
assign R_LUT[124]=14'b00011011110010;
assign R_LUT[125]=14'b00011101100001;
assign R_LUT[126]=14'b00011111010011;
assign R_LUT[127]=14'b00100001000110;
assign R_LUT[128]=14'b00010000000000;
assign R_LUT[129]=14'b00010000000111;
assign R_LUT[130]=14'b00010000011111;
assign R_LUT[131]=14'b00010001000101;
assign R_LUT[132]=14'b00010001111000;
assign R_LUT[133]=14'b00010010110111;
assign R_LUT[134]=14'b00010100000000;
assign R_LUT[135]=14'b00010101010000;
assign R_LUT[136]=14'b00010110101000;
assign R_LUT[137]=14'b00011000000101;
assign R_LUT[138]=14'b00011001100111;
assign R_LUT[139]=14'b00011011001100;
assign R_LUT[140]=14'b00011100110110;
assign R_LUT[141]=14'b00011110100001;
assign R_LUT[142]=14'b00100000001111;
assign R_LUT[143]=14'b00100010000000;
assign R_LUT[144]=14'b00010010000000;
assign R_LUT[145]=14'b00010010000111;
assign R_LUT[146]=14'b00010010011100;
assign R_LUT[147]=14'b00010010111110;
assign R_LUT[148]=14'b00010011101100;
assign R_LUT[149]=14'b00010100100101;
assign R_LUT[150]=14'b00010101101000;
assign R_LUT[151]=14'b00010110110011;
assign R_LUT[152]=14'b00011000000101;
assign R_LUT[153]=14'b00011001011101;
assign R_LUT[154]=14'b00011010111010;
assign R_LUT[155]=14'b00011100011011;
assign R_LUT[156]=14'b00011110000000;
assign R_LUT[157]=14'b00011111100111;
assign R_LUT[158]=14'b00100001010010;
assign R_LUT[159]=14'b00100010111111;
assign R_LUT[160]=14'b00010100000000;
assign R_LUT[161]=14'b00010100000110;
assign R_LUT[162]=14'b00010100011001;
assign R_LUT[163]=14'b00010100111000;
assign R_LUT[164]=14'b00010101100010;
assign R_LUT[165]=14'b00010110010111;
assign R_LUT[166]=14'b00010111010100;
assign R_LUT[167]=14'b00011000011010;
assign R_LUT[168]=14'b00011001100111;
assign R_LUT[169]=14'b00011010111010;
assign R_LUT[170]=14'b00011100010010;
assign R_LUT[171]=14'b00011101101110;
assign R_LUT[172]=14'b00011111001111;
assign R_LUT[173]=14'b00100000110011;
assign R_LUT[174]=14'b00100010011010;
assign R_LUT[175]=14'b00100100000011;
assign R_LUT[176]=14'b00010110000000;
assign R_LUT[177]=14'b00010110000101;
assign R_LUT[178]=14'b00010110010111;
assign R_LUT[179]=14'b00010110110011;
assign R_LUT[180]=14'b00010111011010;
assign R_LUT[181]=14'b00011000001010;
assign R_LUT[182]=14'b00011001000011;
assign R_LUT[183]=14'b00011010000100;
assign R_LUT[184]=14'b00011011001100;
assign R_LUT[185]=14'b00011100011011;
assign R_LUT[186]=14'b00011101101110;
assign R_LUT[187]=14'b00011111000111;
assign R_LUT[188]=14'b00100000100011;
assign R_LUT[189]=14'b00100010000011;
assign R_LUT[190]=14'b00100011100110;
assign R_LUT[191]=14'b00100101001100;
assign R_LUT[192]=14'b00011000000000;
assign R_LUT[193]=14'b00011000000101;
assign R_LUT[194]=14'b00011000010101;
assign R_LUT[195]=14'b00011000101111;
assign R_LUT[196]=14'b00011001010011;
assign R_LUT[197]=14'b00011010000000;
assign R_LUT[198]=14'b00011010110101;
assign R_LUT[199]=14'b00011011110010;
assign R_LUT[200]=14'b00011100110110;
assign R_LUT[201]=14'b00011110000000;
assign R_LUT[202]=14'b00011111001111;
assign R_LUT[203]=14'b00100000100011;
assign R_LUT[204]=14'b00100001111100;
assign R_LUT[205]=14'b00100011011000;
assign R_LUT[206]=14'b00100100111000;
assign R_LUT[207]=14'b00100110011010;
assign R_LUT[208]=14'b00011010000000;
assign R_LUT[209]=14'b00011010000100;
assign R_LUT[210]=14'b00011010010011;
assign R_LUT[211]=14'b00011010101011;
assign R_LUT[212]=14'b00011011001100;
assign R_LUT[213]=14'b00011011110110;
assign R_LUT[214]=14'b00011100101000;
assign R_LUT[215]=14'b00011101100001;
assign R_LUT[216]=14'b00011110100001;
assign R_LUT[217]=14'b00011111100111;
assign R_LUT[218]=14'b00100000110011;
assign R_LUT[219]=14'b00100010000011;
assign R_LUT[220]=14'b00100011011000;
assign R_LUT[221]=14'b00100100110001;
assign R_LUT[222]=14'b00100110001101;
assign R_LUT[223]=14'b00100111101100;
assign R_LUT[224]=14'b00011100000000;
assign R_LUT[225]=14'b00011100000100;
assign R_LUT[226]=14'b00011100010010;
assign R_LUT[227]=14'b00011100101000;
assign R_LUT[228]=14'b00011101000111;
assign R_LUT[229]=14'b00011101101110;
assign R_LUT[230]=14'b00011110011101;
assign R_LUT[231]=14'b00011111010011;
assign R_LUT[232]=14'b00100000001111;
assign R_LUT[233]=14'b00100001010010;
assign R_LUT[234]=14'b00100010011010;
assign R_LUT[235]=14'b00100011100110;
assign R_LUT[236]=14'b00100100111000;
assign R_LUT[237]=14'b00100110001101;
assign R_LUT[238]=14'b00100111100110;
assign R_LUT[239]=14'b00101001000010;
assign R_LUT[240]=14'b00011110000000;
assign R_LUT[241]=14'b00011110000100;
assign R_LUT[242]=14'b00011110010000;
assign R_LUT[243]=14'b00011110100110;
assign R_LUT[244]=14'b00011111000011;
assign R_LUT[245]=14'b00011111100111;
assign R_LUT[246]=14'b00100000010011;
assign R_LUT[247]=14'b00100001000110;
assign R_LUT[248]=14'b00100010000000;
assign R_LUT[249]=14'b00100010111111;
assign R_LUT[250]=14'b00100100000011;
assign R_LUT[251]=14'b00100101001100;
assign R_LUT[252]=14'b00100110011010;
assign R_LUT[253]=14'b00100111101100;
assign R_LUT[254]=14'b00101001000010;
assign R_LUT[255]=14'b00101010011011;

/*****************************************************************/
// Adder Look up table 
assign adder_LUT[0]=4'b0010;
assign adder_LUT[1]=4'b0010;
assign adder_LUT[2]=4'b0011;
assign adder_LUT[3]=4'b0010;
assign adder_LUT[4]=4'b0011;
assign adder_LUT[5]=4'b0011;
assign adder_LUT[6]=4'b0100;
assign adder_LUT[7]=4'b0010;
assign adder_LUT[8]=4'b0011;
assign adder_LUT[9]=4'b0011;
assign adder_LUT[10]=4'b0100;
assign adder_LUT[11]=4'b0011;
assign adder_LUT[12]=4'b0100;
assign adder_LUT[13]=4'b0100;
assign adder_LUT[14]=4'b0101;
assign adder_LUT[15]=4'b0010;
assign adder_LUT[16]=4'b0010;
assign adder_LUT[17]=4'b0010;
assign adder_LUT[18]=4'b0011;
assign adder_LUT[19]=4'b0010;
assign adder_LUT[20]=4'b0011;
assign adder_LUT[21]=4'b0011;
assign adder_LUT[22]=4'b0100;
assign adder_LUT[23]=4'b0010;
assign adder_LUT[24]=4'b0011;
assign adder_LUT[25]=4'b0011;
assign adder_LUT[26]=4'b0100;
assign adder_LUT[27]=4'b011;
assign adder_LUT[28]=4'b0100;
assign adder_LUT[29]=4'b0100;
assign adder_LUT[30]=4'b0101;
assign adder_LUT[31]=4'b0010;
assign adder_LUT[32]=4'b0011;
assign adder_LUT[33]=4'b0011;
assign adder_LUT[34]=4'b0100;
assign adder_LUT[35]=4'b0011;
assign adder_LUT[36]=4'b0100;
assign adder_LUT[37]=4'b0100;
assign adder_LUT[38]=4'b0101;
assign adder_LUT[39]=4'b0011;
assign adder_LUT[40]=4'b0100;
assign adder_LUT[41]=4'b0100;
assign adder_LUT[42]=4'b0101;
assign adder_LUT[43]=4'b0100;
assign adder_LUT[44]=4'b0101;
assign adder_LUT[45]=4'b0101;
assign adder_LUT[46]=4'b0110;
assign adder_LUT[47]=4'b0011;
assign adder_LUT[48]=4'b0010;
assign adder_LUT[49]=4'b0010;
assign adder_LUT[50]=4'b0011;
assign adder_LUT[51]=4'b0010;
assign adder_LUT[52]=4'b0011;
assign adder_LUT[53]=4'b0011;
assign adder_LUT[54]=4'b0100;
assign adder_LUT[55]=4'b0010;
assign adder_LUT[56]=4'b0011;
assign adder_LUT[57]=4'b0011;
assign adder_LUT[58]=4'b0100;
assign adder_LUT[59]=4'b0011;
assign adder_LUT[60]=4'b0100;
assign adder_LUT[61]=4'b0100;
assign adder_LUT[62]=4'b0101;
assign adder_LUT[63]=4'b0010;
assign adder_LUT[64]=4'b0011;
assign adder_LUT[65]=4'b0011;
assign adder_LUT[66]=4'b0100;
assign adder_LUT[67]=4'b0011;
assign adder_LUT[68]=4'b0100;
assign adder_LUT[69]=4'b0100;
assign adder_LUT[70]=4'b0101;
assign adder_LUT[71]=4'b0011;
assign adder_LUT[72]=4'b0100;
assign adder_LUT[73]=4'b0100;
assign adder_LUT[74]=4'b0101;
assign adder_LUT[75]=4'b0100;
assign adder_LUT[76]=4'b0101;
assign adder_LUT[77]=4'b0101;
assign adder_LUT[78]=4'b0110;
assign adder_LUT[79]=4'b0011;
assign adder_LUT[80]=4'b0011;
assign adder_LUT[81]=4'b0011;
assign adder_LUT[82]=4'b0100;
assign adder_LUT[83]=4'b0011;
assign adder_LUT[84]=4'b0100;
assign adder_LUT[85]=4'b0100;
assign adder_LUT[86]=4'b0101;
assign adder_LUT[87]=4'b0011;
assign adder_LUT[88]=4'b0100;
assign adder_LUT[89]=4'b0100;
assign adder_LUT[90]=4'b0101;
assign adder_LUT[91]=4'b0100;
assign adder_LUT[92]=4'b0101;
assign adder_LUT[93]=4'b0101;
assign adder_LUT[94]=4'b0110;
assign adder_LUT[95]=4'b0011;
assign adder_LUT[96]=4'b0100;
assign adder_LUT[97]=4'b0100;
assign adder_LUT[98]=4'b0101;
assign adder_LUT[99]=4'b0100;
assign adder_LUT[100]=4'b0101;
assign adder_LUT[101]=4'b0101;
assign adder_LUT[102]=4'b0110;
assign adder_LUT[103]=4'b0100;
assign adder_LUT[104]=4'b0101;
assign adder_LUT[105]=4'b0101;
assign adder_LUT[106]=4'b0110;
assign adder_LUT[107]=4'b0101;
assign adder_LUT[108]=4'b0110;
assign adder_LUT[109]=4'b0110;
assign adder_LUT[110]=4'b0111;
assign adder_LUT[111]=4'b0100;
assign adder_LUT[112]=4'b0010;
assign adder_LUT[113]=4'b0010;
assign adder_LUT[114]=4'b0011;
assign adder_LUT[115]=4'b0010;
assign adder_LUT[116]=4'b0011;
assign adder_LUT[117]=4'b0011;
assign adder_LUT[118]=4'b0100;
assign adder_LUT[119]=4'b0010;
assign adder_LUT[120]=4'b0011;
assign adder_LUT[121]=4'b0011;
assign adder_LUT[122]=4'b0100;
assign adder_LUT[123]=4'b0011;
assign adder_LUT[124]=4'b0100;
assign adder_LUT[125]=4'b0100;
assign adder_LUT[126]=4'b0101;
assign adder_LUT[127]=4'b0010;
assign adder_LUT[128]=4'b0011;
assign adder_LUT[129]=4'b0011;
assign adder_LUT[130]=4'b0100;
assign adder_LUT[131]=4'b0011;
assign adder_LUT[132]=4'b0100;
assign adder_LUT[133]=4'b0100;
assign adder_LUT[134]=4'b0101;
assign adder_LUT[135]=4'b0011;
assign adder_LUT[136]=4'b0100;
assign adder_LUT[137]=4'b0100;
assign adder_LUT[138]=4'b0101;
assign adder_LUT[139]=4'b0100;
assign adder_LUT[140]=4'b0101;
assign adder_LUT[141]=4'b0101;
assign adder_LUT[142]=4'b0110;
assign adder_LUT[143]=4'b0011;
assign adder_LUT[144]=4'b0011;
assign adder_LUT[145]=4'b0011;
assign adder_LUT[146]=4'b0100;
assign adder_LUT[147]=4'b0011;
assign adder_LUT[148]=4'b0100;
assign adder_LUT[149]=4'b0100;
assign adder_LUT[150]=4'b0101;
assign adder_LUT[151]=4'b0011;
assign adder_LUT[152]=4'b0100;
assign adder_LUT[153]=4'b0100;
assign adder_LUT[154]=4'b0101;
assign adder_LUT[155]=4'b0100;
assign adder_LUT[156]=4'b0101;
assign adder_LUT[157]=4'b0101;
assign adder_LUT[158]=4'b0110;
assign adder_LUT[159]=4'b0011;
assign adder_LUT[160]=4'b0100;
assign adder_LUT[161]=4'b0100;
assign adder_LUT[162]=4'b0101;
assign adder_LUT[163]=4'b0100;
assign adder_LUT[164]=4'b0101;
assign adder_LUT[165]=4'b0101;
assign adder_LUT[166]=4'b0110;
assign adder_LUT[167]=4'b0100;
assign adder_LUT[168]=4'b0101;
assign adder_LUT[169]=4'b0101;
assign adder_LUT[170]=4'b0110;
assign adder_LUT[171]=4'b0101;
assign adder_LUT[172]=4'b0110;
assign adder_LUT[173]=4'b0110;
assign adder_LUT[174]=4'b0111;
assign adder_LUT[175]=4'b0100;
assign adder_LUT[176]=4'b0011;
assign adder_LUT[177]=4'b0011;
assign adder_LUT[178]=4'b0100;
assign adder_LUT[179]=4'b0011;
assign adder_LUT[180]=4'b0100;
assign adder_LUT[181]=4'b0100;
assign adder_LUT[182]=4'b0101;
assign adder_LUT[183]=4'b0011;
assign adder_LUT[184]=4'b0100;
assign adder_LUT[185]=4'b0100;
assign adder_LUT[186]=4'b0101;
assign adder_LUT[187]=4'b0100;
assign adder_LUT[188]=4'b0101;
assign adder_LUT[189]=4'b0101;
assign adder_LUT[190]=4'b0110;
assign adder_LUT[191]=4'b0011;
assign adder_LUT[192]=4'b0100;
assign adder_LUT[193]=4'b0100;
assign adder_LUT[194]=4'b0101;
assign adder_LUT[195]=4'b0100;
assign adder_LUT[196]=4'b0101;
assign adder_LUT[197]=4'b0101;
assign adder_LUT[198]=4'b0110;
assign adder_LUT[199]=4'b0100;
assign adder_LUT[200]=4'b0101;
assign adder_LUT[201]=4'b0101;
assign adder_LUT[202]=4'b0110;
assign adder_LUT[203]=4'b0101;
assign adder_LUT[204]=4'b0110;
assign adder_LUT[205]=4'b0110;
assign adder_LUT[206]=4'b0111;
assign adder_LUT[207]=4'b0100;
assign adder_LUT[208]=4'b0100;
assign adder_LUT[209]=4'b0100;
assign adder_LUT[210]=4'b0101;
assign adder_LUT[211]=4'b0100;
assign adder_LUT[212]=4'b0101;
assign adder_LUT[213]=4'b0101;
assign adder_LUT[214]=4'b0110;
assign adder_LUT[215]=4'b0100;
assign adder_LUT[216]=4'b0101;
assign adder_LUT[217]=4'b0101;
assign adder_LUT[218]=4'b0110;
assign adder_LUT[219]=4'b0101;
assign adder_LUT[220]=4'b0110;
assign adder_LUT[221]=4'b0110;
assign adder_LUT[222]=4'b0111;
assign adder_LUT[223]=4'b0100;
assign adder_LUT[224]=4'b0101;
assign adder_LUT[225]=4'b0101;
assign adder_LUT[226]=4'b0110;
assign adder_LUT[227]=4'b0101;
assign adder_LUT[228]=4'b0110;
assign adder_LUT[229]=4'b0110;
assign adder_LUT[230]=4'b0111;
assign adder_LUT[231]=4'b0101;
assign adder_LUT[232]=4'b0110;
assign adder_LUT[233]=4'b0110;
assign adder_LUT[234]=4'b0111;
assign adder_LUT[235]=4'b0110;
assign adder_LUT[236]=4'b0111;
assign adder_LUT[237]=4'b0111;
assign adder_LUT[238]=4'b1000;
assign adder_LUT[239]=4'b0101;
assign adder_LUT[240]=4'b0010;
assign adder_LUT[241]=4'b0010;
assign adder_LUT[242]=4'b00011;
assign adder_LUT[243]=4'b0010;
assign adder_LUT[244]=4'b0011;
assign adder_LUT[245]=4'b0011;
assign adder_LUT[246]=4'b0100;
assign adder_LUT[247]=4'b0010;
assign adder_LUT[248]=4'b0011;
assign adder_LUT[249]=4'b0011;
assign adder_LUT[250]=4'b0100;
assign adder_LUT[251]=4'b0011;
assign adder_LUT[252]=4'b0100;
assign adder_LUT[253]=4'b0100;
assign adder_LUT[254]=4'b0101;
assign adder_LUT[255]=4'b0010;

/*******************************************************/	
// Tan Look up table	 
assign tan_LUT[0]=14'b10110100000000;
assign tan_LUT[1]=14'b10110100000000;
assign tan_LUT[2]=14'b10110100000000;
assign tan_LUT[3]=14'b10110100000000;
assign tan_LUT[4]=14'b10110100000000;
assign tan_LUT[5]=14'b10110100000000;
assign tan_LUT[6]=14'b10110100000000;
assign tan_LUT[7]=14'b10110100000000;
assign tan_LUT[8]=14'b10110100000000;
assign tan_LUT[9]=14'b10110100000000;
assign tan_LUT[10]=14'b10110100000000;
assign tan_LUT[11]=14'b10110100000000;
assign tan_LUT[12]=14'b10110100000000;
assign tan_LUT[13]=14'b10110100000000;
assign tan_LUT[14]=14'b10110100000000;
assign tan_LUT[15]=14'b10110100000000;
assign tan_LUT[16]=14'b00000000000000;
assign tan_LUT[17]=14'b01011010000000;
assign tan_LUT[18]=14'b01111110110111;
assign tan_LUT[19]=14'b10001111001000;
assign tan_LUT[20]=14'b10010111111011;
assign tan_LUT[21]=14'b10011101011000;
assign tan_LUT[22]=14'b10100001000100;
assign tan_LUT[23]=14'b10100011101111;
assign tan_LUT[24]=14'b10100101110000;
assign tan_LUT[25]=14'b10100111010100;
assign tan_LUT[26]=14'b10101000100101;
assign tan_LUT[27]=14'b10101001100111;
assign tan_LUT[28]=14'b10101010011110;
assign tan_LUT[29]=14'b10101011001100;
assign tan_LUT[30]=14'b10101011110101;
assign tan_LUT[31]=14'b10101100010111;
assign tan_LUT[32]=14'b00000000000000;
assign tan_LUT[33]=14'b00110101001000;
assign tan_LUT[34]=14'b01011010000000;
assign tan_LUT[35]=14'b01110000100111;
assign tan_LUT[36]=14'b01111110110111;
assign tan_LUT[37]=14'b10001000011001;
assign tan_LUT[38]=14'b10001111001000;
assign tan_LUT[39]=14'b10010100000110;
assign tan_LUT[40]=14'b10010111111011;
assign tan_LUT[41]=14'b10011010111100;
assign tan_LUT[42]=14'b10011101011000;
assign tan_LUT[43]=14'b10011111011000;
assign tan_LUT[44]=14'b10100001000100;
assign tan_LUT[45]=14'b10100010100000;
assign tan_LUT[46]=14'b10100011101111;
assign tan_LUT[47]=14'b10100100110011;
assign tan_LUT[48]=14'b00000000000000;
assign tan_LUT[49]=14'b00100100110111;
assign tan_LUT[50]=14'b01000011011000;
assign tan_LUT[51]=14'b01011010000000;
assign tan_LUT[52]=14'b01101010010000;
assign tan_LUT[53]=14'b01110110000100;
assign tan_LUT[54]=14'b01111110110111;
assign tan_LUT[55]=14'b10000101100110;
assign tan_LUT[56]=14'b10001010111000;
assign tan_LUT[57]=14'b10001111001000;
assign tan_LUT[58]=14'b10010010100110;
assign tan_LUT[59]=14'b10010101011111;
assign tan_LUT[60]=14'b10010111111011;
assign tan_LUT[61]=14'b10011010000000;
assign tan_LUT[62]=14'b10011011110011;
assign tan_LUT[63]=14'b10011101011000;
assign tan_LUT[64]=14'b00000000000000;
assign tan_LUT[65]=14'b00011100000100;
assign tan_LUT[66]=14'b00110101001000;
assign tan_LUT[67]=14'b01001001101111;
assign tan_LUT[68]=14'b01011010000000;
assign tan_LUT[69]=14'b01100110101011;
assign tan_LUT[70]=14'b01110000100111;
assign tan_LUT[71]=14'b01111000100000;
assign tan_LUT[72]=14'b01111110110111;
assign tan_LUT[73]=14'b10000100000100;
assign tan_LUT[74]=14'b10001000011001;
assign tan_LUT[75]=14'b10001100000010;
assign tan_LUT[76]=14'b10001111001000;
assign tan_LUT[77]=14'b10010001110010;
assign tan_LUT[78]=14'b10010100000110;
assign tan_LUT[79]=14'b10010110001000;
assign tan_LUT[80]=14'b00000000000000;
assign tan_LUT[81]=14'b00010110100111;
assign tan_LUT[82]=14'b00101011100110;
assign tan_LUT[83]=14'b00111101111011;
assign tan_LUT[84]=14'b01001101010100;
assign tan_LUT[85]=14'b01011010000000;
assign tan_LUT[86]=14'b01100100011000;
assign tan_LUT[87]=14'b01101100111011;
assign tan_LUT[88]=14'b01110011111111;
assign tan_LUT[89]=14'b01111001111001;
assign tan_LUT[90]=14'b01111110110111;
assign tan_LUT[91]=14'b10000011000111;
assign tan_LUT[92]=14'b10000110110000;
assign tan_LUT[93]=14'b10001001111011;
assign tan_LUT[94]=14'b10001100101100;
assign tan_LUT[95]=14'b10001111001000;
assign tan_LUT[96]=14'b00000000000000;
assign tan_LUT[97]=14'b00010010111011;
assign tan_LUT[98]=14'b00100100110111;
assign tan_LUT[99]=14'b00110101001000;
assign tan_LUT[100]=14'b01000011011000;
assign tan_LUT[101]=14'b01001111100111;
assign tan_LUT[102]=14'b01011010000000;
assign tan_LUT[103]=14'b01100010110011;
assign tan_LUT[104]=14'b01101010010000;
assign tan_LUT[105]=14'b01110000100111;
assign tan_LUT[106]=14'b01110110000100;
assign tan_LUT[107]=14'b01111010110001;
assign tan_LUT[108]=14'b01111110110111;
assign tan_LUT[109]=14'b10000010011100;
assign tan_LUT[110]=14'b10000101100110;
assign tan_LUT[111]=14'b10001000011001;
assign tan_LUT[112]=14'b00000000000000;
assign tan_LUT[113]=14'b00010000010000;
assign tan_LUT[114]=14'b00011111111001;
assign tan_LUT[115]=14'b00101110011001;
assign tan_LUT[116]=14'b00111011011111;
assign tan_LUT[117]=14'b01000111000100;
assign tan_LUT[118]=14'b01010001001100;
assign tan_LUT[119]=14'b01011010000000;
assign tan_LUT[120]=14'b01100001101000;
assign tan_LUT[121]=14'b01101000010000;
assign tan_LUT[122]=14'b01101110000001;
assign tan_LUT[123]=14'b01110011000011;
assign tan_LUT[124]=14'b01110111011111;
assign tan_LUT[125]=14'b01111011011001;
assign tan_LUT[126]=14'b01111110110111;
assign tan_LUT[127]=14'b10000001111101;
assign tan_LUT[128]=14'b00000000000000;
assign tan_LUT[129]=14'b00001110010000;
assign tan_LUT[130]=14'b00011100000100;
assign tan_LUT[131]=14'b00101001000111;
assign tan_LUT[132]=14'b00110101001000;
assign tan_LUT[133]=14'b01000000000000;
assign tan_LUT[134]=14'b01001001101111;
assign tan_LUT[135]=14'b01010010010111;
assign tan_LUT[136]=14'b01011010000000;
assign tan_LUT[137]=14'b01100000101110;
assign tan_LUT[138]=14'b01100110101011;
assign tan_LUT[139]=14'b01101011111100;
assign tan_LUT[140]=14'b01110000100111;
assign tan_LUT[141]=14'b01110100110010;
assign tan_LUT[142]=14'b01111000100000;
assign tan_LUT[143]=14'b01111011110110;
assign tan_LUT[144]=14'b00000000000000;
assign tan_LUT[145]=14'b00001100101011;
assign tan_LUT[146]=14'b00011001000011;
assign tan_LUT[147]=14'b00100100110111;
assign tan_LUT[148]=14'b00101111111011;
assign tan_LUT[149]=14'b00111010000110;
assign tan_LUT[150]=14'b01000011011000;
assign tan_LUT[151]=14'b01001011110000;
assign tan_LUT[152]=14'b01010011010001;
assign tan_LUT[153]=14'b01011010000000;
assign tan_LUT[154]=14'b01100000000001;
assign tan_LUT[155]=14'b01100101011010;
assign tan_LUT[156]=14'b01101010010000;
assign tan_LUT[157]=14'b01101110100111;
assign tan_LUT[158]=14'b01110010100001;
assign tan_LUT[159]=14'b01110110000100;
assign tan_LUT[160]=14'b00000000000000;
assign tan_LUT[161]=14'b00001011011010;
assign tan_LUT[162]=14'b00010110100111;
assign tan_LUT[163]=14'b00100001011001;
assign tan_LUT[164]=14'b00101011100110;
assign tan_LUT[165]=14'b00110101001000;
assign tan_LUT[166]=14'b00111101111011;
assign tan_LUT[167]=14'b01000101111110;
assign tan_LUT[168]=14'b01001101010100;
assign tan_LUT[169]=14'b01010011111110;
assign tan_LUT[170]=14'b01011010000000;
assign tan_LUT[171]=14'b01011111011100;
assign tan_LUT[172]=14'b01100100011000;
assign tan_LUT[173]=14'b01101000110111;
assign tan_LUT[174]=14'b01101100111011;
assign tan_LUT[175]=14'b01110000100111;
assign tan_LUT[176]=14'b00000000000000;
assign tan_LUT[177]=14'b00001010011000;
assign tan_LUT[178]=14'b00010100100111;
assign tan_LUT[179]=14'b00011110100000;
assign tan_LUT[180]=14'b00100111111101;
assign tan_LUT[181]=14'b00110000111000;
assign tan_LUT[182]=14'b00111001001110;
assign tan_LUT[183]=14'b01000000111100;
assign tan_LUT[184]=14'b01001000000011;
assign tan_LUT[185]=14'b01001110100101;
assign tan_LUT[186]=14'b01010100100011;
assign tan_LUT[187]=14'b01011010000000;
assign tan_LUT[188]=14'b01011110111110;
assign tan_LUT[189]=14'b01100011100001;
assign tan_LUT[190]=14'b01100111101011;
assign tan_LUT[191]=14'b01101011011111;
assign tan_LUT[192]=14'b00000000000000;
assign tan_LUT[193]=14'b00001001100001;
assign tan_LUT[194]=14'b00010010111011;
assign tan_LUT[195]=14'b00011100000100;
assign tan_LUT[196]=14'b00100100110111;
assign tan_LUT[197]=14'b00101101001111;
assign tan_LUT[198]=14'b00110101001000;
assign tan_LUT[199]=14'b00111100100000;
assign tan_LUT[200]=14'b01000011011000;
assign tan_LUT[201]=14'b01001001101111;
assign tan_LUT[202]=14'b01001111100111;
assign tan_LUT[203]=14'b01010101000001;
assign tan_LUT[204]=14'b01011010000000;
assign tan_LUT[205]=14'b01011110100101;
assign tan_LUT[206]=14'b01100010110011;
assign tan_LUT[207]=14'b01100110101011;
assign tan_LUT[208]=14'b00000000000000;
assign tan_LUT[209]=14'b00001000110011;
assign tan_LUT[210]=14'b00010001011111;
assign tan_LUT[211]=14'b00011001111111;
assign tan_LUT[212]=14'b00100010001101;
assign tan_LUT[213]=14'b00101010000100;
assign tan_LUT[214]=14'b00110001100011;
assign tan_LUT[215]=14'b00111000100110;
assign tan_LUT[216]=14'b00111111001101;
assign tan_LUT[217]=14'b01000101011000;
assign tan_LUT[218]=14'b01001011001000;
assign tan_LUT[219]=14'b01010000011110;
assign tan_LUT[220]=14'b01010101011010;
assign tan_LUT[221]=14'b01011010000000;
assign tan_LUT[222]=14'b01011110001111;
assign tan_LUT[223]=14'b01100010001010;
assign tan_LUT[224]=14'b00000000000000;
assign tan_LUT[225]=14'b00001000001010;
assign tan_LUT[226]=14'b00010000010000;
assign tan_LUT[227]=14'b00011000001100;
assign tan_LUT[228]=14'b00011111111001;
assign tan_LUT[229]=14'b00100111010011;
assign tan_LUT[230]=14'b00101110011001;
assign tan_LUT[231]=14'b00110101001000;
assign tan_LUT[232]=14'b00111011011111;
assign tan_LUT[233]=14'b01000001011110;
assign tan_LUT[234]=14'b01000111000100;
assign tan_LUT[235]=14'b01001100010100;
assign tan_LUT[236]=14'b01010001001100;
assign tan_LUT[237]=14'b01010101110000;
assign tan_LUT[238]=14'b01011010000000;
assign tan_LUT[239]=14'b01011101111100;
assign tan_LUT[240]=14'b00000000000000;
assign tan_LUT[241]=14'b00000111101000;
assign tan_LUT[242]=14'b00001111001100;
assign tan_LUT[243]=14'b00010110100111;
assign tan_LUT[244]=14'b00011101110111;
assign tan_LUT[245]=14'b00100100110111;
assign tan_LUT[246]=14'b00101011100110;
assign tan_LUT[247]=14'b00110010000010;
assign tan_LUT[248]=14'b00111000001001;
assign tan_LUT[249]=14'b00111101111011;
assign tan_LUT[250]=14'b01000011011000;
assign tan_LUT[251]=14'b01001000100000;
assign tan_LUT[252]=14'b01001101010100;
assign tan_LUT[253]=14'b01010001110101;
assign tan_LUT[254]=14'b01010110000011;
assign tan_LUT[255]=14'b01011010000000;

/************************************************/
//Define Inputs and Outputs
input clk;
input [13:0] R_fixed ;
input [13:0] angle1;
input [13:0] angle2;
input [3:0] adder;
input [4:0] error;
output [7:0] final_cord1 ;
output [7:0] final_cord2 ;

/************************************************/
//Define other temporary variables 	
reg [13:0] data_outR; 
reg [13:0] data_outtan; 
reg [3:0] data_outadder; 
reg [7:0] count=8'b00000000;
reg [9:0] globalcount=9'b000000000;
reg [3:0] count1=4'b0000;
reg [3:0] globalcount1=4'b0000;
reg [13:0] deltaAngle1=14'b00000000000000;
reg [13:0] deltaAngle2=14'b00000000000000;
reg [14:0] deltaAdd=15'b000000000000000;
reg [14:0] AngleMin=15'b111111111111111;
reg [13:0] temp = 14'b00000000000000;
reg [13:0] temp1 = 14'b00000000000000;
reg [3:0] flag1=4'b0000;
reg [3:0] flag2=4'b0000;
reg [7:0] counter_1 [9:0] ;
reg [13:0] counter_R_1 [9:0] ;
reg [7:0] counter_2 [9:0] ;
reg [13:0] counter_R_2 [9:0] ;
reg [7:0] final_cord1=8'b00000000;
reg [7:0] final_cord2=8'b00000000;
reg [13:0] subtract_R = 14'b11111111111111;
reg [3:0] X = 4'b0000;
reg [3:0] Y = 4'b0000;
reg [3:0] X1 = 4'b0000;
reg [3:0] Y1 = 4'b0000;
reg [7:0] final_count_1 = 8'b00000000;
reg [7:0] final_count_2 = 8'b00000000;

/*****************************************************************/
// Clock triggered always block
always@(posedge clk)
begin
	//If globalcount value is less than 764 
	if(globalcount < 764)
	begin
		//Increment globalcount
		globalcount=globalcount+1;
		//Sequential block is triggered after every 4th clock cycle 
		if(globalcount==1 || globalcount==4 || globalcount==7 || globalcount==10 || globalcount==13 || globalcount==16 || globalcount==19 || globalcount==22 || globalcount==25 || globalcount==28 || globalcount==31 || globalcount==34 || globalcount==37 || globalcount==40 || globalcount==43 || globalcount==46 || globalcount==49 || globalcount==52 || globalcount==55 || globalcount==58 || globalcount==61 || globalcount==64 || globalcount==67 || globalcount==70 || globalcount==73 || globalcount==76 || globalcount==79 || globalcount==82 || globalcount==85 || globalcount==88 || globalcount==91 || globalcount==94 || globalcount==97 ||globalcount==100 || globalcount==103 || globalcount==106 || globalcount==109 || globalcount==112 || globalcount==115 || globalcount==118 || globalcount==121 || globalcount==124 || globalcount==127 || globalcount==130 || globalcount==133 || globalcount==136 || globalcount==139 || globalcount==142 || globalcount==145 || globalcount==148 || globalcount==151 || globalcount==154 || globalcount==157 || globalcount==160 || globalcount==163 || globalcount==166 || globalcount==169 || globalcount==172 || globalcount==175 || globalcount==178 || globalcount==181 || globalcount==184 || globalcount==187 || globalcount==190 || globalcount==193 || globalcount==196 || globalcount==199 || globalcount==202 || globalcount==205 || globalcount==208 || globalcount==211 || globalcount==214 || globalcount==217 || globalcount==220 || globalcount==223 || globalcount==226 || globalcount==229 || globalcount==232 || globalcount==235 || globalcount==238 || globalcount==241 || globalcount==244 || globalcount==247 || globalcount==250 || globalcount==253 || globalcount==256 || globalcount==259 || globalcount==262 || globalcount==265 || globalcount==268 || globalcount==271 || globalcount==274 || globalcount==277 || globalcount==280 || globalcount==283 || globalcount==286 || globalcount==289 || globalcount==292 || globalcount==295 || globalcount==298 || globalcount==301 || globalcount==304 || globalcount==307 || globalcount==310 || globalcount==313 || globalcount==316 || globalcount==319 || globalcount==322 || globalcount==325 || globalcount==328 || globalcount==331 || globalcount==334 || globalcount==337 || globalcount==340 || globalcount==343 || globalcount==346 || globalcount==349 || globalcount==352 || globalcount==355 || globalcount==358 || globalcount==361 || globalcount==364 || globalcount==367 || globalcount==370 || globalcount==373 || globalcount==376 || globalcount==379 || globalcount==382 || globalcount==385 || globalcount==388 || globalcount==391 || globalcount==394 || globalcount==397 || globalcount==400 || globalcount==403 || globalcount==406 || globalcount==409 || globalcount==412 || globalcount==415 || globalcount==418 || globalcount==421 || globalcount==424 || globalcount==427 || globalcount==430 || globalcount==433 || globalcount==436 || globalcount==439 || globalcount==442 || globalcount==445 || globalcount==448 || globalcount==451 || globalcount==454 || globalcount==457 || globalcount==460 || globalcount==463 ||globalcount==466 || globalcount==469 || globalcount==472 || globalcount==475 || globalcount==478 || globalcount==481 || globalcount==484 || globalcount==487 || globalcount==490 || globalcount==493 || globalcount==496 || globalcount==499 || globalcount==502 || globalcount==505 || globalcount==508 || globalcount==511 || globalcount==514 || globalcount==517 || globalcount==520 || globalcount==523 || globalcount==526 || globalcount==529 || globalcount==532 || globalcount==535 || globalcount==538 || globalcount==541 || globalcount==544 || globalcount==547 || globalcount==550 || globalcount==553 || globalcount==556 || globalcount==559 || globalcount==562 || globalcount==565 || globalcount==568 || globalcount==571 || globalcount==574 || globalcount==577 || globalcount==580 || globalcount==583 || globalcount==586 || globalcount==589 || globalcount==592 || globalcount==595 || globalcount==598 || globalcount==601 || globalcount==604 || globalcount==607 || globalcount==610 || globalcount==613 || globalcount==616 || globalcount==619 || globalcount==622 || globalcount==625 || globalcount==628 || globalcount==631 || globalcount==634 || globalcount==637 || globalcount==640 || globalcount==643 || globalcount==646 || globalcount==649 || globalcount==652 || globalcount==655 || globalcount==658 || globalcount==661 || globalcount==664 || globalcount==667 || globalcount==670 || globalcount==673 || globalcount==676 || globalcount==679 || globalcount==682 || globalcount==685 || globalcount==688 || globalcount==691 || globalcount==694 || globalcount==697 || globalcount==700 || globalcount==703 || globalcount==706 || globalcount==709 || globalcount==712 || globalcount==715 || globalcount==718 || globalcount==721 || globalcount==724 || globalcount==727 || globalcount==730 ||globalcount==733 ||globalcount==736 || globalcount==739 || globalcount==742 || globalcount==745 || globalcount==748 || globalcount==751 || globalcount==754 || globalcount==757 || globalcount==760 || globalcount==763) 
		begin
			count = count + 8'b00000001;
			//Read data from memory i.e. R value from R_LUT, tan value from tan_LUT and adder value from adder_LUT
			data_outR = R_LUT[count];
			data_outadder = adder_LUT[count];
			data_outtan = tan_LUT[count];
			//Taking positive difference of data_outtan and angle1
			temp=(data_outtan>angle1)?(data_outtan-angle1):(angle1-data_outtan);
			//Checking for conditions of values of R, tan and adders to find a few near to optimum coordinates for angle1
			if(data_outR < R_fixed  && data_outadder < adder && (temp)< sind_LUT[error])
			begin
				//Storing values of count and R for each value which satisfies the above conditions
				counter_1[flag1]=count;
				counter_R_1[flag1]=data_outR;
				flag1=flag1+4'b0001;
			end

			//Taking positive difference of data_outtan and angle2
			temp1=(data_outtan>angle2)?(data_outtan-angle2):(angle2-data_outtan);
			//Checking for conditions of values of R, tan and adders to find a few near to optimum coordinates for angle2
			if(data_outR < R_fixed  && data_outadder < adder && (temp1)< sind_LUT[error])
			begin
				//Storing values of count and R for each value which satisfies the above conditions
				counter_2[flag2]=count;
				counter_R_2[flag2]=data_outR;
				flag2=flag2+4'b0001;
			end
		end
	end
	//After all possible values of coordinates have been accessed we get 2 arrays one per angle with a few near to optimum coordinate values. Else will then find the optimum most point for the same
	else 
	begin
	 if(globalcount1 != flag1)
	 begin
		//Taking positive difference of R's of both the angles written to the memory in previous step
		temp1=(counter_R_2[globalcount1]>counter_R_1[count1])?(counter_R_2[globalcount1]-counter_R_1[count1]):(counter_R_1[count1]-counter_R_2[globalcount1]);
		//Find the coordinates one for each angle such as the difference between their absolutes values i.e. R values is the minimum. Also for points having same value of difference of their absolute value a point with least angular error is selected
		if(temp1 < subtract_R)
		begin
			subtract_R =temp1;
			final_count_1 = counter_1[globalcount1];
			final_count_2 = counter_2[count1];
			deltaAngle1=tan_LUT[final_count_1]-angle1;
			deltaAngle2=tan_LUT[final_count_2]-angle2;
			deltaAdd=deltaAngle1+deltaAngle2;
			if(deltaAdd<AngleMin)
			begin
				AngleMin=deltaAdd;
				final_cord1=counter_1[globalcount1];
				final_cord2=counter_2[count1];
			end
			count1=count1+4'b0001;
			
		end
		if(count1==flag2)
		begin
			count1=0;
			globalcount1=globalcount1+4'b0001;
		end
	 end	
	end
end
endmodule
